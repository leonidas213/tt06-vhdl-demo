LIBRARY IEEE;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity controllogic is
  port (
    a      : in  std_logic;
    b      : in  std_logic;
    c      : in  std_logic;
    d      : in  std_logic;
    e      : in  std_logic;
    f      : in  std_logic;
    g      : in  std_logic;
    muxb0  : out std_logic;
    muxb1  : out std_logic;
    muxb2  : out std_logic;
    src2d  : out std_logic;
    aluop0 : out std_logic;
    aluop1 : out std_logic;
    aluop2 : out std_logic;
    aluop3 : out std_logic;
    aluop4 : out std_logic;
    we     : out std_logic;
    sf     : out std_logic;
    alu2d  : out std_logic;
    iem0   : out std_logic;
    iem1   : out std_logic;
    br0    : out std_logic;
    br1    : out std_logic;
    br2    : out std_logic;
    muxa   : out std_logic;
    ld     : out std_logic;
    st     : out std_logic;
    p_abs  : out std_logic;
    iow    : out std_logic;
    ior    : out std_logic;
    stpc   : out std_logic;
    reti   : out std_logic;
    rand   : out std_logic);
end entity;

architecture behavioral of controllogic is
  signal s0 : std_logic;
  signal s1 : std_logic;
  signal s2 : std_logic;
  signal s3 : std_logic;
  signal s4 : std_logic;
  signal s5 : std_logic;
  signal s6 : std_logic;
begin
  s5     <= not a;
  s0     <= not b;
  s1     <= not c;
  s2     <= not d;
  s3     <= not e;
  s6     <= not f;
  s4     <= not g;
  muxb0  <= ((a and s0 and s1 and s2 and s3 and f and s4) or (a and s0 and s1 and s2 and e and f and g) or (s5 and s1 and d and e and f and s4) or (s5 and b and c and s3 and s6 and s4) or (s5 and s0 and s1 and d and f and s4) or (s5 and s0 and s1 and d and e and s4) or (s5 and s0 and c and s2 and s3 and s4) or (s5 and b and s1 and s2 and s3 and g) or (s5 and c and d and s6 and g) or (s5 and c and s2 and e and g) or (s5 and b and c and e and g) or (s5 and b and c and s2 and e));
  muxb1  <= ((a and s0 and s1 and s2 and e and f and s4) or (s5 and c and s2 and s3 and s6 and g) or (s5 and b and s1 and s2 and s3 and s4) or (a and s0 and s1 and s2 and s3 and g) or (a and s0 and s1 and s2 and s3 and s6) or (s5 and s1 and d and f and g) or (s5 and c and d and s6 and s4) or (s5 and b and c and s6 and g) or (s5 and b and c and f and s4) or (s5 and c and s2 and e and s4) or (s5 and s0 and s1 and d and g) or (s5 and b and d and e) or (s5 and b and c and e));
  muxb2  <= ((s5 and b and c and d and e and f and g) or (s5 and c and s2 and s3 and s6 and s4) or (s5 and b and s2 and s3 and f and g) or (s5 and b and s1 and s3 and f and g) or (s5 and s0 and s1 and d and f and s4) or (s5 and s0 and c and d and s6 and g) or (a and s0 and s1 and s2 and f and g) or (s5 and s0 and c and s2 and s3 and s4) or (s5 and s0 and c and s2 and e and g) or (s5 and b and s1 and s2 and s3 and g) or (a and s0 and s1 and s2 and s3 and s4) or (s5 and s1 and d and e and s4));
  src2d  <= ((s5 and s0 and s1 and s2 and s3 and s6 and g) or (s5 and b and s1 and d and s3 and f and g) or (s5 and b and s1 and d and e and s6 and g) or (s5 and b and c and s2 and s3 and s6 and g) or (a and s0 and s1 and s2 and s3 and s6 and s4) or (s5 and b and d and e and f and s4) or (s5 and b and c and d and e and f));
  aluop0 <= ((s5 and s0 and s1 and d and e and f and s4) or (s5 and s0 and c and s2 and s3 and s6 and g) or (s5 and s0 and c and s2 and s3 and f and s4) or (s5 and s0 and c and d and e and f and g) or (s5 and s1 and s2 and s3 and f and g) or (s5 and s0 and s1 and e and s6 and g) or (s5 and b and s1 and s2 and f));
  aluop1 <= ((s5 and s0 and c and d and s3 and f and g) or (a and s0 and s1 and s2 and e and s6 and g) or (a and s0 and s1 and s2 and e and f and s4) or (s5 and b and s1 and d and s3 and s4) or (s5 and s0 and c and d and e and s6) or (s5 and b and s1 and d and s3 and s6) or (s5 and b and s1 and s2 and e));
  aluop2 <= ((s5 and b and s1 and d and s3 and f and s4) or (a and s0 and s1 and s2 and e and s6 and g) or (a and s0 and s1 and s2 and e and f and s4) or (s5 and s0 and s2 and e and f and g) or (s5 and s0 and d and s3 and s6 and s4) or (s5 and s0 and c and s3 and f and g) or (s5 and s0 and c and s2 and e and f) or (s5 and s0 and c and d and s6) or (s5 and s0 and c and d and s3));
  aluop3 <= ((s5 and s0 and d and e and f and g) or (s5 and s0 and c and d and f and s4) or (s5 and s0 and s2 and e and s6) or (s5 and b and s1 and s3 and s6) or (s5 and s0 and c and s2 and s3) or (s5 and b and s1 and s2 and s3) or (s0 and s1 and s2 and e and s6 and g) or (s0 and s1 and s2 and e and f and s4));
  aluop4 <= ((s5 and b and c and s2 and s3 and s6 and g) or (s5 and b and c and s2 and s3 and f and s4) or (a and s0 and s1 and s2 and s3 and s6 and s4) or (s5 and s1 and d and e and s6 and s4) or (s5 and s0 and s1 and e and f and s4) or (s5 and s0 and s1 and s2 and f and s4) or (s5 and s0 and c and d and s3 and g) or (s5 and b and s1 and s2 and e and g) or (s5 and b and s1 and d and s3 and g) or (s5 and s0 and s3 and f and g) or (s5 and s0 and d and s6 and s4) or (s5 and s0 and d and e and s6) or (s5 and s0 and c and e and s6) or (s0 and s1 and s2 and s3 and f and g));
  we     <= ((s5 and d and s3 and f and s4) or (s5 and s1 and e and s6 and s4) or (s5 and s1 and e and f and g) or (s5 and c and s2 and s3 and s4) or (s5 and s1 and d and s3 and s6) or (s5 and c and s2 and s3 and f) or (s5 and s0 and d and s6) or (s5 and s1 and s2 and e) or (s5 and s0 and d and s3) or (s5 and s0 and s1 and d) or (s5 and s0 and c and s2) or (s0 and s1 and s2 and g) or (s0 and s1 and s2 and f));
  sf     <= ((s5 and s1 and d and s3 and s6 and s4) or (s5 and s0 and s2 and f and s4) or (s5 and s0 and d and f and g) or (s5 and s0 and s1 and f and g) or (s5 and s0 and c and s6) or (s5 and b and s1 and s2) or (s5 and s0 and e) or (s0 and s1 and s2 and e and s6 and g) or (s0 and s1 and s2 and e and f and s4));
  alu2d  <= ((s5 and c and s2 and s3 and f and g) or (s5 and s1 and d and s3 and s4) or (s5 and s1 and d and s3 and s6) or (s5 and s0 and e and s6) or (s5 and s0 and s2 and f) or (s5 and s0 and s1 and f) or (s5 and s1 and s2 and e) or (s5 and s0 and c and s3) or (s0 and s1 and s2 and e and s6 and g) or (s0 and s1 and s2 and e and f and s4));
  iem0   <= ((s5 and s0 and c and s2 and s3 and s6 and g) or (a and s0 and s1 and s2 and s3 and s6 and g) or (a and s0 and s1 and s2 and e and f and s4) or (s5 and c and d and e and s6 and s4) or (s5 and s0 and c and d and s6 and s4) or (s5 and b and c and d and f and s4) or (s5 and s0 and c and s2 and e and s4) or (s5 and b and s1 and s2 and s3 and s4) or (s5 and s1 and d and e and g) or (s5 and s0 and s1 and d and g));
  iem1   <= ((s5 and b and s1 and d and e and s6 and g) or (s5 and b and c and d and e and f and s4));
  br0    <= ((s5 and b and c and s2 and e and f and g) or (s5 and b and c and d and s6 and g) or (s5 and b and c and d and s3 and s6));
  br1    <= ((s5 and b and c and s2 and e and s6 and g) or (s5 and b and c and s2 and e and f and s4) or (s5 and b and c and d and s3 and s6));
  br2    <= ((s5 and b and c and d and s3 and s6 and g) or (s5 and b and c and s2 and e and s4) or (s5 and b and c and s2 and e and f));
  muxa   <= ((s5 and b and s1 and d and e and s6 and s4) or (s5 and b and c and s2 and s3 and f and s4) or (a and s0 and s1 and s2 and s3 and g) or (a and s0 and s1 and s2 and s3 and f));
  ld     <= ((s5 and b and s1 and d and e and s6 and s4) or (s5 and b and s1 and d and e and f and g) or (s5 and b and c and s2 and s3 and s4));
  st     <= ((s5 and b and s1 and d and s3 and f and g) or (s5 and b and s1 and d and e and s6 and g) or (s5 and b and s1 and d and e and f and s4) or (s5 and b and c and s2 and s3 and s6 and g));
  p_abs  <= ((s5 and b and c and d and e and s6 and s4) or (a and s0 and s1 and s2 and e and s6 and s4) or (s5 and b and c and d and s3 and f));
  iow    <= ((a and s0 and s1 and s2 and s3 and s6 and s4) or (s5 and b and c and d and e and f));
  ior    <= ((a and s0 and s1 and s2 and s3 and g) or (a and s0 and s1 and s2 and s3 and f));
  stpc   <= (s5 and b and c and d and s3 and f and s4);
  reti   <= (a and s0 and s1 and s2 and e and s6 and s4);
  rand   <= (a and s0 and s1 and s2 and e and f and g);
end architecture;

